module sumador_4_y_1(  
	input [3:0] in_sum, 
	output [3:0] out_sum 
);
	assign  out_sum=in_sum+1;
endmodule